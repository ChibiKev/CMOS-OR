*** SPICE deck for cell 2-input_NOR{lay} from library Project1
*** Created on Fri Sep 20, 2019 16:20:04
*** Last revised on Fri Sep 20, 2019 17:42:50
*** Written on Fri Sep 20, 2019 17:43:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: 2-input_NOR{lay}
Mnmos@0 gnd A Vout gnd NMOS L=0.35U W=1.75U AS=1.48P AD=4.364P PS=4.025U PD=12.075U
Mnmos@1 Vout B gnd gnd NMOS L=0.35U W=1.75U AS=4.364P AD=1.48P PS=12.075U PD=4.025U
Mpmos@0 vdd A net@0 vdd PMOS L=0.35U W=1.75U AS=1.914P AD=6.738P PS=3.937U PD=18.375U
Mpmos@1 net@0 B Vout vdd PMOS L=0.35U W=1.75U AS=1.48P AD=1.914P PS=4.025U PD=3.937U

* Spice Code nodes in cell cell '2-input_NOR{lay}'
VDD VDD 0 DC 3.3
VGND GND 0 DC 0
Vin A 0 PULSE (3.3 0 0 0.01n 0.01n 10n 20n)
Vin2 B 0 PULSE (3.3 0 0 0.01n 0.01n 20n 40n)
.TRAN 0 50n
.include C:\Users\kille\Desktop\Electric\C5_models.txt
.END
